CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 D:\Online Classes\CircuitMaker2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
52
13 Logic Switch~
5 746 522 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5433 0 0
2
5.89968e-315 0
0
13 Logic Switch~
5 691 132 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3679 0 0
2
5.89968e-315 5.26354e-315
0
13 Logic Switch~
5 109 536 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9342 0 0
2
44201.5 0
0
13 Logic Switch~
5 111 490 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3623 0 0
2
44201.5 1
0
13 Logic Switch~
5 112 406 0 1 11
0 42
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3722 0 0
2
44201.5 2
0
13 Logic Switch~
5 110 368 0 1 11
0 43
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8993 0 0
2
44201.5 3
0
13 Logic Switch~
5 112 300 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3723 0 0
2
44201.5 4
0
13 Logic Switch~
5 113 253 0 1 11
0 45
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6244 0 0
2
44201.5 5
0
13 Logic Switch~
5 110 150 0 1 11
0 46
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6421 0 0
2
44201.5 6
0
13 Logic Switch~
5 110 103 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7743 0 0
2
44201.5 7
0
8 3-In OR~
219 596 528 0 4 22
0 3 4 5 2
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
9840 0 0
2
44201.5 8
0
14 Logic Display~
6 1112 504 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6910 0 0
2
5.89968e-315 5.30499e-315
0
14 Logic Display~
6 1110 438 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
449 0 0
2
5.89968e-315 5.32571e-315
0
8 2-In OR~
219 987 524 0 3 22
0 8 7 48
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 10 0
1 U
8761 0 0
2
5.89968e-315 5.34643e-315
0
9 2-In AND~
219 921 514 0 3 22
0 9 10 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
6748 0 0
2
5.89968e-315 5.3568e-315
0
6 74136~
219 911 456 0 3 22
0 10 9 6
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
7393 0 0
2
5.89968e-315 5.36716e-315
0
9 2-In AND~
219 813 506 0 3 22
0 12 11 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
7699 0 0
2
5.89968e-315 5.37752e-315
0
6 74136~
219 809 447 0 3 22
0 11 12 10
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
6638 0 0
2
5.89968e-315 5.38788e-315
0
14 Logic Display~
6 1117 296 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
5.89968e-315 5.39306e-315
0
8 2-In OR~
219 1003 391 0 3 22
0 15 14 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
9395 0 0
2
5.89968e-315 5.39824e-315
0
9 2-In AND~
219 936 382 0 3 22
0 17 16 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3303 0 0
2
5.89968e-315 5.40342e-315
0
6 74136~
219 928 328 0 3 22
0 16 17 13
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U8D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
4498 0 0
2
5.89968e-315 5.4086e-315
0
9 2-In AND~
219 815 393 0 3 22
0 18 2 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
9728 0 0
2
5.89968e-315 5.41378e-315
0
6 74136~
219 807 341 0 3 22
0 2 18 17
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U8C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3789 0 0
2
5.89968e-315 5.41896e-315
0
8 2-In OR~
219 999 250 0 3 22
0 20 19 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3978 0 0
2
5.89968e-315 5.42414e-315
0
14 Logic Display~
6 1053 158 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3494 0 0
2
5.89968e-315 5.42933e-315
0
9 2-In AND~
219 941 241 0 3 22
0 23 22 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3507 0 0
2
5.89968e-315 5.43192e-315
0
6 74136~
219 935 188 0 3 22
0 22 23 21
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U8B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
5151 0 0
2
5.89968e-315 5.43451e-315
0
14 Logic Display~
6 1057 47 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
5.89968e-315 5.4371e-315
0
9 2-In AND~
219 786 249 0 3 22
0 25 2 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
8585 0 0
2
5.89968e-315 5.43969e-315
0
6 74136~
219 779 198 0 3 22
0 25 2 23
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U8A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
8809 0 0
2
5.89968e-315 5.44228e-315
0
9 2-In AND~
219 863 138 0 3 22
0 26 27 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
5993 0 0
2
44201.5 9
0
6 74136~
219 853 87 0 3 22
0 27 26 24
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8654 0 0
2
44201.5 10
0
9 2-In AND~
219 547 417 0 3 22
0 25 12 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7223 0 0
2
44201.5 11
0
9 2-In AND~
219 485 478 0 3 22
0 18 12 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3641 0 0
2
44201.5 12
0
8 2-In OR~
219 386 536 0 3 22
0 29 28 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3104 0 0
2
44201.5 13
0
9 2-In AND~
219 321 526 0 3 22
0 30 31 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3296 0 0
2
44201.5 14
0
6 74136~
219 312 488 0 3 22
0 31 30 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8534 0 0
2
44201.5 15
0
8 2-In OR~
219 381 414 0 3 22
0 33 32 30
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
949 0 0
2
44201.5 16
0
9 2-In AND~
219 322 406 0 3 22
0 35 34 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3371 0 0
2
44201.5 17
0
6 74136~
219 317 366 0 3 22
0 35 34 18
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7311 0 0
2
44201.5 18
0
8 2-In OR~
219 382 294 0 3 22
0 37 36 34
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3409 0 0
2
44201.5 19
0
9 2-In AND~
219 329 284 0 3 22
0 38 39 37
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3526 0 0
2
44201.5 20
0
6 74136~
219 322 244 0 3 22
0 38 39 25
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4129 0 0
2
44201.5 21
0
6 74136~
219 207 481 0 3 22
0 40 41 31
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6278 0 0
2
44201.5 22
0
9 2-In AND~
219 206 545 0 3 22
0 40 41 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3482 0 0
2
44201.5 23
0
9 2-In AND~
219 220 415 0 3 22
0 42 43 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8323 0 0
2
44201.5 24
0
6 74136~
219 216 358 0 3 22
0 43 42 35
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3984 0 0
2
44201.5 25
0
9 2-In AND~
219 220 307 0 3 22
0 45 44 36
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7622 0 0
2
44201.5 26
0
6 74136~
219 216 242 0 3 22
0 45 44 39
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
816 0 0
2
44201.5 27
0
9 2-In AND~
219 224 156 0 3 22
0 47 46 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4656 0 0
2
44201.5 28
0
6 74136~
219 221 86 0 3 22
0 47 46 27
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6356 0 0
2
44201.5 29
0
80
1 0 2 0 0 8320 0 12 0 0 5 4
1112 522
1112 598
708 598
708 524
2 0 2 0 0 0 0 23 0 0 5 2
791 402
708 402
1 0 2 0 0 0 0 24 0 0 5 2
791 332
708 332
2 0 2 0 0 0 0 30 0 0 5 2
762 258
708 258
4 2 2 0 0 128 0 11 31 0 0 4
629 528
708 528
708 207
763 207
3 1 3 0 0 8320 0 34 11 0 0 4
568 417
579 417
579 519
583 519
3 2 4 0 0 12416 0 35 11 0 0 4
506 478
524 478
524 528
584 528
3 3 5 0 0 8320 0 36 11 0 0 3
419 536
419 537
583 537
3 1 6 0 0 4224 0 16 13 0 0 2
944 456
1110 456
3 2 7 0 0 8320 0 17 14 0 0 3
834 506
834 533
974 533
3 1 8 0 0 8320 0 15 14 0 0 3
942 514
942 515
974 515
0 1 9 0 0 4096 0 0 15 13 0 3
883 465
883 505
897 505
3 2 9 0 0 12416 0 20 16 0 0 6
1036 391
1066 391
1066 416
883 416
883 465
895 465
0 2 10 0 0 4224 0 0 15 15 0 3
867 447
867 523
897 523
3 1 10 0 0 0 0 18 16 0 0 2
842 447
895 447
0 1 11 0 0 4224 0 0 18 17 0 3
783 515
783 438
793 438
1 2 11 0 0 0 0 1 17 0 0 4
758 522
783 522
783 515
789 515
0 1 12 0 0 4096 0 0 17 19 0 3
761 456
761 497
789 497
0 2 12 0 0 8320 0 0 18 44 0 3
511 426
511 456
793 456
3 1 13 0 0 4224 0 22 19 0 0 3
961 328
1117 328
1117 314
3 2 14 0 0 12416 0 23 20 0 0 4
836 393
856 393
856 400
990 400
3 1 15 0 0 4224 0 21 20 0 0 2
957 382
990 382
1 0 16 0 0 4096 0 22 0 0 24 2
912 319
881 319
3 2 16 0 0 12416 0 25 21 0 0 6
1032 250
1055 250
1055 296
881 296
881 391
912 391
0 1 17 0 0 4096 0 0 21 26 0 3
902 341
902 373
912 373
3 2 17 0 0 4224 0 24 22 0 0 4
840 341
903 341
903 337
912 337
0 1 18 0 0 8192 0 0 23 28 0 3
761 366
761 384
791 384
0 2 18 0 0 4224 0 0 24 45 0 4
459 366
761 366
761 350
791 350
3 2 19 0 0 8320 0 30 25 0 0 3
807 249
807 259
986 259
3 1 20 0 0 4224 0 27 25 0 0 2
962 241
986 241
3 1 21 0 0 4224 0 28 26 0 0 3
968 188
1053 188
1053 176
0 2 22 0 0 4224 0 0 27 33 0 3
900 179
900 250
917 250
3 1 22 0 0 0 0 32 28 0 0 4
884 138
900 138
900 179
919 179
0 1 23 0 0 8192 0 0 27 35 0 3
851 197
851 232
917 232
3 2 23 0 0 8320 0 31 28 0 0 3
812 198
812 197
919 197
3 1 24 0 0 4224 0 33 29 0 0 3
886 87
1057 87
1057 65
0 1 25 0 0 4096 0 0 30 38 0 3
506 244
762 244
762 240
0 1 25 0 0 8320 0 0 31 43 0 3
506 244
506 189
763 189
0 1 26 0 0 4096 0 0 32 40 0 3
825 132
839 132
839 129
1 2 26 0 0 4224 0 2 33 0 0 4
703 132
827 132
827 96
837 96
0 2 27 0 0 8192 0 0 32 42 0 3
737 78
737 147
839 147
3 1 27 0 0 4224 0 52 33 0 0 4
254 86
725 86
725 78
837 78
3 1 25 0 0 0 0 44 34 0 0 4
355 244
509 244
509 408
523 408
0 2 12 0 0 0 0 0 34 46 0 3
455 487
455 426
523 426
3 1 18 0 0 0 0 41 35 0 0 3
350 366
461 366
461 469
3 2 12 0 0 0 0 38 35 0 0 3
345 488
345 487
461 487
3 2 28 0 0 4224 0 46 36 0 0 2
227 545
373 545
3 1 29 0 0 8320 0 37 36 0 0 3
342 526
342 527
373 527
0 1 30 0 0 8192 0 0 37 50 0 3
276 497
276 517
297 517
3 2 30 0 0 12416 0 39 38 0 0 6
414 414
447 414
447 458
276 458
276 497
296 497
0 2 31 0 0 4224 0 0 37 52 0 3
247 479
247 535
297 535
3 1 31 0 0 0 0 45 38 0 0 3
240 481
240 479
296 479
3 2 32 0 0 12416 0 47 39 0 0 4
241 415
254 415
254 423
368 423
3 1 33 0 0 8320 0 40 39 0 0 3
343 406
343 405
368 405
0 2 34 0 0 4096 0 0 40 56 0 3
277 373
277 415
298 415
3 2 34 0 0 12416 0 42 41 0 0 6
415 294
442 294
442 325
277 325
277 375
301 375
0 1 35 0 0 8192 0 0 40 58 0 3
255 357
255 397
298 397
3 1 35 0 0 8320 0 48 41 0 0 3
249 358
249 357
301 357
3 2 36 0 0 4224 0 49 42 0 0 4
241 307
359 307
359 303
369 303
3 1 37 0 0 8320 0 43 42 0 0 3
350 284
350 285
369 285
0 1 38 0 0 4096 0 0 43 62 0 3
292 235
292 275
305 275
3 1 38 0 0 8320 0 51 44 0 0 4
245 156
292 156
292 235
306 235
0 2 39 0 0 4224 0 0 43 64 0 3
268 251
268 293
305 293
3 2 39 0 0 0 0 50 44 0 0 4
249 242
268 242
268 253
306 253
0 1 40 0 0 4224 0 0 45 66 0 3
160 536
160 472
191 472
1 1 40 0 0 0 0 3 46 0 0 2
121 536
182 536
0 2 41 0 0 4096 0 0 46 68 0 3
137 490
137 554
182 554
1 2 41 0 0 4224 0 4 45 0 0 2
123 490
191 490
0 2 42 0 0 4096 0 0 48 70 0 3
178 406
178 367
200 367
1 1 42 0 0 4224 0 5 47 0 0 2
124 406
196 406
0 2 43 0 0 8320 0 0 47 72 0 3
133 368
133 424
196 424
1 1 43 0 0 0 0 6 48 0 0 4
122 368
147 368
147 349
200 349
0 2 44 0 0 4224 0 0 50 75 0 3
164 316
164 251
200 251
0 1 45 0 0 4224 0 0 49 76 0 3
186 233
186 298
196 298
1 2 44 0 0 0 0 7 49 0 0 4
124 300
148 300
148 316
196 316
1 1 45 0 0 0 0 8 50 0 0 4
125 253
148 253
148 233
200 233
0 2 46 0 0 4224 0 0 52 79 0 3
175 165
175 95
205 95
0 1 47 0 0 8192 0 0 51 80 0 3
147 103
147 147
200 147
1 2 46 0 0 0 0 9 51 0 0 4
122 150
140 150
140 165
200 165
1 1 47 0 0 12416 0 10 52 0 0 4
122 103
148 103
148 77
205 77
28
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
677 544 706 568
687 552 695 568
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
357 334 394 358
367 342 383 358
2 Z4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
341 454 378 478
351 462 367 478
2 Z8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
424 386 461 410
434 394 450 410
2 C3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
407 547 436 571
417 555 425 571
1 K
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
349 198 386 222
359 206 375 222
2 Z2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
417 259 454 283
427 267 443 283
2 C2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
273 37 310 61
283 45 299 61
2 Z1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
253 121 290 145
263 129 279 145
2 C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
62 522 99 546
72 530 88 546
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
57 464 94 488
67 472 83 488
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
59 397 96 421
69 405 85 421
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
62 351 99 375
72 359 88 375
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
59 281 96 305
69 289 85 305
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
58 228 95 252
68 236 84 252
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
52 125 89 149
62 133 78 149
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
47 76 84 100
57 84 73 100
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
642 118 671 142
652 126 660 142
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1087 40 1124 64
1097 48 1113 64
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1098 147 1135 171
1108 155 1124 171
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1161 276 1198 300
1171 284 1187 300
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
920 111 965 135
930 119 954 135
3 C1'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1049 219 1094 243
1059 227 1083 243
3 C2'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
949 335 994 359
959 343 983 359
3 C3'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
732 527 761 551
742 535 750 551
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1136 416 1173 440
1146 424 1162 440
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1142 498 1187 522
1152 506 1176 522
3 C4'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
433 607 710 631
443 615 699 631
32 BCD Adder with basic logic gates
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
